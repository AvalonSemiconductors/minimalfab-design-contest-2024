* Created by KLayout

* cell TOP
.SUBCKT TOP
* device instance $1 r0 *1 371,32 PMOS
M$1 28 7 22 22 PMOS L=10U W=30U AS=570P AD=570P PS=98U PD=98U
* device instance $2 r0 *1 183,32 PMOS
M$2 29 6 23 23 PMOS L=10U W=30U AS=570P AD=375P PS=98U PD=55U
* device instance $3 r0 *1 218,32 PMOS
M$3 27 5 29 29 PMOS L=10U W=30U AS=375P AD=570P PS=55U PD=98U
* device instance $4 r0 *1 277,32 PMOS
M$4 30 4 25 25 PMOS L=10U W=30U AS=570P AD=375P PS=98U PD=55U
* device instance $5 r0 *1 312,32 PMOS
M$5 31 3 30 30 PMOS L=10U W=30U AS=375P AD=570P PS=55U PD=98U
* device instance $6 r0 *1 124,32 PMOS
M$6 32 3 26 26 PMOS L=10U W=30U AS=570P AD=570P PS=98U PD=98U
* device instance $7 r0 *1 24,32 PMOS
M$7 21 1 24 24 PMOS L=10U W=30U AS=570P AD=450P PS=98U PD=60U
* device instance $8 r0 *1 64,32 PMOS
M$8 33 2 21 21 PMOS L=10U W=30U AS=450P AD=570P PS=60U PD=98U
* device instance $9 r0 *1 277,-66.5 NMOS
M$9 19 4 13 13 NMOS L=10U W=10U AS=190P AD=125P PS=58U PD=35U
* device instance $10 r0 *1 312,-66.5 NMOS
M$10 20 5 19 19 NMOS L=10U W=10U AS=125P AD=190P PS=35U PD=58U
* device instance $11 r0 *1 371,-66.5 NMOS
M$11 18 7 12 12 NMOS L=10U W=10U AS=190P AD=190P PS=58U PD=58U
* device instance $12 r0 *1 24,-66.5 NMOS
M$12 8 1 9 9 NMOS L=10U W=10U AS=190P AD=150P PS=58U PD=40U
* device instance $13 r0 *1 64,-66.5 NMOS
M$13 14 2 8 8 NMOS L=10U W=10U AS=150P AD=190P PS=40U PD=58U
* device instance $14 r0 *1 183,-66.5 NMOS
M$14 16 6 11 11 NMOS L=10U W=10U AS=190P AD=125P PS=58U PD=35U
* device instance $15 r0 *1 218,-66.5 NMOS
M$15 17 3 16 16 NMOS L=10U W=10U AS=125P AD=190P PS=35U PD=58U
* device instance $16 r0 *1 124,-66.5 NMOS
M$16 15 3 10 10 NMOS L=10U W=10U AS=190P AD=190P PS=58U PD=58U
.ENDS TOP
